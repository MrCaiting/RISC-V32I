import rv32i_types::*;

module cache_control
(

    );

endmodule : cache_control
