library verilog;
use verilog.vl_types.all;
entity write_cache_sv_unit is
end write_cache_sv_unit;
